training@here.6171
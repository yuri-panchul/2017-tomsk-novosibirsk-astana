`ifdef word_width
`else
`define word_width 16
`endif

`ifdef stack_size
`else
`define stack_size 4
`endif

`ifdef stack_pointer_size
`else
`define stack_pointer_size 2
`endif
